`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:32:25 08/05/2021 
// Design Name: 
// Module Name:    E 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module E(
    input [31:0] E_instr,
    input [31:0] E_PC,
    input [31:0] E_RS_DATA,
    input [31:0] E_RT_DATA,
    input [31:0] E_EXTDATA
    );

    

endmodule
